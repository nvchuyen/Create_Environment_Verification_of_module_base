
//---------------------------------------
//
//---------------------------------------
`ifndef DFF_IF
`define DFF_IF

interface dff_if;
  logic clk;
  logic rst;
  logic din;
  logic dout;
endinterface : dff_if

`endif
